THERMO
  300.   1000.   4000.
HE                      HE  1               G    300.00   4000.00 1000.00      1
 .250000000E+01 .000000000E+00 .000000000E+00 .000000000E+00 .000000000E+00    2
-.745375000E+03 .928723974E+00 .250000000E+01 .000000000E+00 .000000000E+00    3
 .000000000E+00 .000000000E+00-.745375000E+03 .928723974E+00                   4
AR                      AR  1               G    300.00   4000.00 1000.00      1
 .250000000E+01 .000000000E+00 .000000000E+00 .000000000E+00 .000000000E+00    2
-.745375000E+03 .436600000E+01 .250000000E+01 .000000000E+00 .000000000E+00    3
 .000000000E+00 .000000000E+00-.745375000E+03 .436600000E+01                   4
N2                      N   2               G    300.00   4000.00 1000.00      1
 .292663788E+01 .148797700E-02-.568476030E-06 .100970400E-09-.675335090E-14    2
-.922795384E+03 .598054018E+01 .329867700E+01 .140823990E-02-.396322180E-05    3
 .564151480E-08-.244485400E-11-.102090000E+04 .395037200E+01                   4
NO                      O   1N   1          G    300.00   4000.00 1000.00      1
 .324543589E+01 .126913800E-02-.501589000E-06 .916928270E-10-.627541890E-14    2
 .980084032E+04 .641728767E+01 .337654100E+01 .125306300E-02-.330275000E-05    3
 .521781020E-08-.244626190E-11 .981796100E+04 .582959200E+01                   4
N2O                     O   1N   2          G    300.00   4000.00 1000.00      1
 .471897567E+01 .287371290E-02-.119749600E-05 .225055100E-09-.157533690E-13    2
 .816581343E+04-.165723704E+01 .254305700E+01 .949219330E-02-.979277500E-05    3
 .626384410E-08-.190182510E-11 .876510200E+04 .951122400E+01                   4
O2                      O   2               G    300.00   4000.00 1000.00      1
 .369757685E+01 .613519690E-03-.125884200E-06 .177528100E-10-.113643500E-14    2
-.123392966E+04 .318917125E+01 .321293600E+01 .112748610E-02-.575614990E-06    3
 .131387700E-08-.876855390E-12-.100524900E+04 .603473900E+01                   4
NO2                     O   2N   1          G    300.00   4000.00 1000.00      1
 .468285677E+01 .246242900E-02-.104225900E-05 .197690200E-09-.139171700E-13    2
 .226129300E+04 .988610659E+00 .267060000E+01 .783849970E-02-.806386380E-05    3
 .616171380E-08-.232014990E-11 .289629000E+04 .116120700E+02                   4
HNO                     H   1O   1N   1     G    300.00   4000.00 1000.00      1
 .361514436E+01 .321248500E-02-.126033690E-05 .226729700E-09-.153623600E-13    2
 .106619122E+05 .481025325E+01 .278440200E+01 .660964610E-02-.930022270E-05    3
 .943798020E-08-.375314580E-11 .109187800E+05 .903562900E+01                   4
HNNO                    H   1O   1N   2     G    300.00   4000.00 1500.00      1
 .699121930E+01 .187597000E-02-.212458400E-06-.671047200E-10 .123050800E-13    2
 .249756641E+05-.112352384E+02 .223829800E+01 .135920000E-01-.117987300E-04    3
 .539297100E-08-.101085900E-11 .266025900E+05 .141367900E+02                   4
HONO                    H   1O   2N   1     G    300.00   4000.00 1000.00      1
 .548688978E+01 .421806500E-02-.164914300E-05 .297187700E-09-.202114800E-13    2
-.112686489E+05-.299698546E+01 .229041300E+01 .140992200E-01-.136787200E-04    3
 .749878000E-08-.187690500E-11-.104319500E+05 .132807700E+02                   4
HNO2                    H   1O   2N   1     G    300.00   4000.00 1500.00      1
 .647962840E+01 .199527400E-02-.174038700E-06-.969587200E-10 .170148000E-13    2
-.999926943E+04-.106728455E+02 .193483800E+01 .101003600E-01-.496461600E-05    3
 .870112000E-09-.232413500E-14-.810548400E+04 .147325000E+02                   4
HONO2                   H   1O   3N   1     G    300.00   4000.00 1500.00      1
 .975613289E+01 .190094800E-02-.324002000E-06-.397663900E-10 .110033400E-13    2
-.194224157E+05-.269001236E+02 .787766800E+00 .238232900E-01-.220596400E-04    3
 .103404800E-07-.197285700E-11-.163044200E+05 .210896400E+02                   4
H2                      H   2               G    300.00   4000.00 1000.00      1
 .299142220E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033546E+03-.135510641E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
N2H2                    H   2N   2          G    300.00   4000.00 1000.00      1
 .337118994E+01 .603996800E-02-.230385300E-05 .406278900E-09-.271314400E-13    2
 .241817095E+05 .498055769E+01 .161799940E+01 .130631220E-01-.171571100E-04    3
 .160560790E-07-.609363800E-11 .246752600E+05 .137946700E+02                   4
H2O                     H   2O   1          G    300.00   4000.00 1000.00      1
 .267214569E+01 .305629290E-02-.873026070E-06 .120099600E-09-.639161790E-14    2
-.298992115E+05 .686281125E+01 .338684200E+01 .347498200E-02-.635469590E-05    3
 .696858040E-08-.250658800E-11-.302081100E+05 .259023200E+01                   4
H2O2                    H   2O   2          G    300.00   4000.00 1000.00      1
 .457316594E+01 .433613590E-02-.147468900E-05 .234890300E-09-.143165410E-13    2
-.180069531E+05 .501137915E+00 .338875300E+01 .656922580E-02-.148501200E-06    3
-.462580510E-08 .247151410E-11-.176631400E+05 .678536300E+01                   4
NH3                     H   3N   1          G    300.00   4000.00 1000.00      1
 .246189456E+01 .605916650E-02-.200497610E-05 .313600310E-09-.193831700E-13    2
-.649326483E+04 .747215046E+01 .220435100E+01 .101147600E-01-.146526500E-04    3
 .144723500E-07-.532850890E-11-.652548900E+04 .812714000E+01                   4
N2H4                    H   4N   2          G    300.00   4000.00 1000.00      1
 .497732211E+01 .959551900E-02-.354763900E-05 .612429900E-09-.402979500E-13    2
 .934121983E+04-.296302077E+01 .644260600E-01 .274973000E-01-.289945100E-04    3
 .174524000E-07-.442228200E-11 .104519200E+05 .212778900E+02                   4
CO                      C   1O   1          G    300.00   4000.00 1000.00      1
 .302507617E+01 .144268900E-02-.563082720E-06 .101858100E-09-.691095110E-14    2
-.142683499E+05 .610822521E+01 .326245100E+01 .151194100E-02-.388175520E-05    3
 .558194380E-08-.247495100E-11-.143105400E+05 .484889700E+01                   4
CO2                     C   1O   2          G    300.00   4000.00 1000.00      1
 .445362582E+01 .314016800E-02-.127841100E-05 .239399610E-09-.166903300E-13    2
-.489669524E+05-.955420007E+00 .227572400E+01 .992207230E-02-.104091100E-04    3
 .686668590E-08-.211728010E-11-.483731400E+05 .101884900E+02                   4
HCN                     C   1H   1N   1     G    300.00   4000.00 1000.00      1
 .365007798E+01 .346099790E-02-.127427900E-05 .221765490E-09-.147717700E-13    2
 .149839102E+05 .239321426E+01 .249046200E+01 .861127950E-02-.103103400E-04    3
 .748149810E-08-.222910900E-11 .152083400E+05 .790498000E+01                   4
HOCN                    C   1H   1O   1N   1G    300.00   4000.00 1000.00      1
 .564560836E+01 .229820610E-02-.216262900E-06-.121480100E-09 .223863610E-13    2
-.317811025E+04-.359027798E+01 .362829200E+01 .566418420E-02-.117020600E-06    3
-.234863800E-08 .801640220E-12-.247592500E+04 .747682300E+01                   4
HCNO                    C   1H   1O   1N   1G    300.00   4000.00 1000.00      1
 .669241213E+01 .236836030E-02-.237151000E-06-.127550300E-09 .240713700E-13    2
 .169473623E+05-.124543537E+02 .318485800E+01 .975231640E-02-.128020300E-05    3
-.616310380E-08 .322627490E-11 .179790700E+05 .612384200E+01                   4
HNCO                    C   1H   1O   1N   1G    300.00   4000.00 1000.00      1
 .621186395E+01 .229713690E-02-.221612790E-06-.122204400E-09 .227240590E-13    2
-.147707257E+05-.801661658E+01 .369405900E+01 .665723530E-02-.505446810E-07    3
-.347341090E-08 .136056900E-11-.139197600E+05 .571273900E+01                   4
CH2O                    C   1H   2O   1     G    300.00   4000.00 1000.00      1
 .299560858E+01 .668132120E-02-.262895400E-05 .473715290E-09-.321251710E-13    2
-.153203666E+05 .691256052E+01 .165273100E+01 .126314400E-01-.188816790E-04    3
 .205003110E-07-.841323710E-11-.148654000E+05 .137848200E+02                   4
HCOOH                   C   1H   2O   2     G    300.00   4000.00 1376.00      1
 .668733013E+01 .514289368E-02-.182238513E-05 .289719163E-09-.170892199E-13    2
-.483995400E+05-.113104798E+02 .143548185E+01 .163363016E-01-.106257421E-04    3
 .332132977E-08-.402176103E-12-.464616504E+05 .172885798E+02                   4
HCO3H                   C   1H   2O   3     G    300.00   4000.00 1378.00      1
 .987503581E+01 .464663708E-02-.167230522E-05 .268624413E-09-.159595232E-13    2
-.380502456E+05-.224938942E+02 .242464726E+01 .219706380E-01-.168705546E-04    3
 .625612194E-08-.911645843E-12-.354828006E+05 .175027796E+02                   4
CH3NO                   C   1H   3O   1N   1G    300.00   4000.00 1500.00      1
 .882055478E+01 .370623300E-02-.289474100E-06-.189791000E-09 .323754400E-13    2
 .536285603E+04-.221322539E+02 .210995500E+01 .151782200E-01-.707178900E-05    3
 .151061100E-08-.160420400E-12 .829361200E+04 .156970200E+02                   4
CH3NO2                  C   1H   3O   2N   1G    300.00   4000.00 1382.00      1
 .673034758E+01 .109601272E-01-.405357875E-05 .667102246E-09-.404686823E-13    2
-.129143475E+05-.101800883E+02 .354053638E+01 .186559899E-02 .444946580E-04    3
-.587057133E-07 .230684496E-10-.111385976E+05 .106884657E+02                   4
CH3ONO                  C   1H   3O   2N   1G    300.00   4000.00 1500.00      1
 .113612738E+02 .415934900E-02-.414567000E-06-.169514000E-09 .302873200E-13    2
-.128147952E+05-.354542296E+02 .149034500E+01 .264543300E-01-.211233200E-04    3
 .941439900E-08-.181120500E-11-.912578200E+04 .181376600E+02                   4
CH3ONO2                 C   1H   3O   3N   1G    300.00   4000.00 1500.00      1
 .143618741E+02 .411224300E-02-.511305200E-06-.149643600E-09 .301215600E-13    2
-.197243835E+05-.513183467E+02 .780335400E+00 .345420400E-01-.282232800E-04    3
 .123232400E-07-.230216400E-11-.146534600E+05 .224575200E+02                   4
CH4                     C   1H   4          G    300.00   4000.00 1000.00      1
 .168346564E+01 .102372400E-01-.387512820E-05 .678558490E-09-.450342310E-13    2
-.100807773E+05 .962347575E+01 .778741700E+00 .174766800E-01-.278340900E-04    3
 .304970800E-07-.122393100E-10-.982522800E+04 .137221900E+02                   4
CH3OH                   C   1H   4O   1     G    300.00   4000.00 1000.00      1
 .402907793E+01 .937659290E-02-.305025380E-05 .435879300E-09-.222472310E-13    2
-.261579223E+05 .237808255E+01 .266011500E+01 .734150780E-02 .717005010E-05    3
-.879319370E-08 .239056990E-11-.253534800E+05 .112326300E+02                   4
CH3OOH                  C   1H   4O   2     G    300.00   4000.00 1000.00      1
 .563694993E+01 .111814780E-01-.369593390E-05 .407189810E-09 .000000000E+00    2
-.180442749E+05-.124166637E+01 .586865100E+01 .107942400E-01-.364552990E-05    3
 .541291180E-09-.289684390E-13-.181268900E+05-.251762300E+01                   4
C2H2                    C   2H   2          G    300.00   4000.00 1000.00      1
 .443677300E+01 .537603910E-02-.191281610E-05 .328637890E-09-.215670900E-13    2
 .256676622E+05-.280035722E+01 .201356200E+01 .151904500E-01-.161631910E-04    3
 .907899180E-08-.191274600E-11 .261244400E+05 .880537800E+01                   4
CH2CO                   C   2H   2O   1     G    300.00   4000.00 1000.00      1
 .603885318E+01 .580484000E-02-.192095400E-05 .279448500E-09-.145886800E-13    2
-.858343402E+04-.765782305E+01 .297497100E+01 .121187100E-01-.234504600E-05    3
-.646668500E-08 .390564900E-11-.763263700E+04 .867355300E+01                   4
C2H2O2                  C   2H   2O   2     G    300.00   4000.00 1386.00      1
 .975438561E+01 .497645947E-02-.174410483E-05 .275586994E-09-.161969892E-13    2
-.295832896E+05-.261878329E+02 .188105120E+01 .236386368E-01-.183443295E-04    3
 .684842963E-08-.992733674E-12-.269280190E+05 .159154793E+02                   4
CH3CN                   C   2H   3N   1     G    300.00   4000.00 1000.00      1
 .239240386E+01 .156188730E-01-.791204970E-05 .193723330E-08-.186119560E-12    2
 .849993803E+04 .111452402E+02 .251975310E+01 .135675230E-01-.257640770E-05    3
-.308939670E-08 .142886920E-11 .855337620E+04 .109208680E+02                   4
C2H4                    C   2H   4          G    300.00   4000.00 1000.00      1
 .352841648E+01 .114851800E-01-.441838480E-05 .784460000E-09-.526684780E-13    2
 .442829030E+04 .223039249E+01-.861487900E+00 .279616190E-01-.338867690E-04    3
 .278515200E-07-.973787890E-11 .557304700E+04 .242114800E+02                   4
C2H4O                   C   2H   4O   1     G    300.00   4000.00 1000.00      1
 .385543260E+01 .146081760E-01-.526121540E-05 .628115500E-09 .000000000E+00    2
-.851874300E+04 .214156911E+01-.130385500E+01 .282461720E-01-.170593430E-04    3
 .394753470E-08 .000000000E+00-.707559900E+04 .289352600E+02                   4
CH3CHO                  C   2H   4O   1     G    300.00   4000.00 1000.00      1
 .586869116E+01 .107942400E-01-.364552990E-05 .541291180E-09-.289684390E-13    2
-.226457128E+05-.601321650E+01 .250569500E+01 .133699100E-01 .467195290E-05    3
-.112814000E-07 .426356610E-11-.212458800E+05 .133508900E+02                   4
C2H4O2                  C   2H   4O   2     G    300.00   4000.00 1358.00      1
 .887306567E+01 .992257253E-02-.334820779E-05 .515546009E-09-.297527820E-13    2
-.410084739E+05-.182786314E+02 .437688685E+01 .159485358E-01-.363672718E-05    3
-.179212805E-08 .741898956E-12-.389689472E+05 .750888268E+01                   4
CH3COOH                 C   2H   4O   2     G    300.00   4000.00 1000.00      1
 .691666936E+01 .128920800E-01-.420990320E-05 .458049540E-09 .000000000E+00    2
-.553508487E+05-.102392103E+02 .846928500E+00 .292145000E-01-.186455200E-04    3
 .464098720E-08 .000000000E+00-.536761800E+05 .211901500E+02                   4
CH3CO3H                 C   2H   4O   3     G    300.00   4000.00 1000.00      1
 .114777196E+02 .831667150E-02-.185084560E-05 .103274160E-09 .000000000E+00    2
-.451075908E+05-.290204723E+02 .484746000E+01 .218580610E-01-.904284660E-05    3
 .384145300E-09 .000000000E+00-.429209100E+05 .674072600E+01                   4
C2-OQOOH                C   2H   4O   3     G    300.00   4000.00 1380.00      1
 .124064339E+02 .947233784E-02-.328107928E-05 .513772211E-09-.299872803E-13    2
-.349123142E+05-.339479874E+02 .552382546E+01 .242068306E-01-.152898974E-04    3
 .501728362E-08-.696406358E-12-.323406789E+05 .357240645E+01                   4
C2H6                    C   2H   6          G    300.00   4000.00 1000.00      1
 .482597579E+01 .138404300E-01-.455725790E-05 .672496720E-09-.359816110E-13    2
-.127178296E+05-.523976258E+01 .146253900E+01 .154946700E-01 .578050690E-05    3
-.125783200E-07 .458626710E-11-.112391800E+05 .144322900E+02                   4
C2H5OH                  C   2H   6O   1     G    300.00   4000.00 1000.00      1
 .434717120E+01 .186288000E-01-.677946700E-05 .816592600E-09 .000000000E+00    2
-.306615743E+05 .324247304E+01 .576535800E+00 .289451200E-01-.161002000E-04    3
 .359164100E-08 .000000000E+00-.296359500E+05 .227081300E+02                   4
C2H5OOH                 C   2H   6O   2     G    300.00   4000.00 1000.00      1
 .914611907E+01 .144611400E-01-.455120020E-05 .475780030E-09 .000000000E+00    2
-.236690607E+05-.205899250E+02 .223998300E+01 .310914290E-01-.170933710E-04    3
 .329379790E-08 .000000000E+00-.216018500E+05 .158174300E+02                   4
C3H2                    C   3H   2          G    300.00   4000.00 1000.00      1
 .767099642E+01 .274874900E-02-.437094300E-06-.645559900E-10 .166388700E-13    2
 .625972092E+05-.123689926E+02 .316671400E+01 .248257200E-01-.459163700E-04    3
 .426801900E-07-.148215200E-10 .635042100E+05 .886944600E+01                   4
AC3H4                   C   3H   4          G    300.00   4000.00 1400.07      1
 .977625145E+01 .530213820E-02-.370111790E-06-.302638610E-09 .508958110E-13    2
 .195497314E+05-.307705909E+02 .253983090E+01 .163343700E-01-.176495000E-05    3
-.464736520E-08 .172913110E-11 .225124300E+05 .993570230E+01                   4
PC3H4                   C   3H   4          G    300.00   4000.00 1000.00      1
 .281460543E+01 .185524496E-01-.955026768E-05 .239951370E-08-.237485257E-12    2
 .207010771E+05 .860604972E+01 .146175323E+01 .246026602E-01-.190219395E-04    3
 .860363422E-08-.166729240E-11 .209209793E+05 .149262585E+02                   4
C2H3CHO                 C   3H   4O   1     G    300.00   4000.00 1393.00      1
 .104184607E+02 .948963321E-02-.329310529E-05 .516279203E-09-.301587291E-13    2
-.149629790E+05-.307232511E+02 .292355162E+00 .354321417E-01-.294936324E-04    3
 .128100124E-07-.226144108E-11-.116521584E+05 .228878280E+02                   4
C3H4O2                  C   3H   4O   2     G    300.00   4000.00 1404.00      1
 .130577477E+02 .906905120E-02-.308189261E-05 .476481380E-09-.275669277E-13    2
-.369274825E+05-.425273740E+02 .147485987E+00 .464706296E-01-.451901760E-04    3
 .219641008E-07-.416219125E-11-.331809255E+05 .242182934E+02                   4
C3H6                    C   3H   6          G    300.00   4000.00 1000.00      1
 .673231663E+01 .149083400E-01-.494989900E-05 .721202210E-09-.376620390E-13    2
-.923623057E+03-.133137684E+02 .149330700E+01 .209251700E-01 .448679380E-05    3
-.166891190E-07 .715814600E-11 .107482600E+04 .161453400E+02                   4
CH3COCH3                C   3H   6O   1     G    300.00   4000.00 1374.00      1
 .991426580E+01 .146030709E-01-.506085765E-05 .792682855E-09-.462739645E-13    2
-.311168055E+05-.286116537E+02 .130767163E+01 .292021742E-01-.119045617E-04    3
 .652150087E-09 .467751203E-12-.275328269E+05 .196395025E+02                   4
C3H6O                   C   3H   6O   1     G    300.00   4000.00 1000.00      1
 .433142310E+01 .236433890E-01-.875060690E-05 .106889830E-08 .000000000E+00    2
-.138496111E+05 .215169726E+01 .507423500E+00 .318789710E-01-.137497700E-04    3
 .165647900E-08 .000000000E+00-.126239100E+05 .226350900E+02                   4
C2H5CHO                 C   3H   6O   1     G    300.00   4000.00 1379.00      1
 .872954858E+01 .199253945E-01-.785642340E-05 .132736406E-08-.812865962E-13    2
-.281462888E+05-.222846545E+02 .441647615E+01 .159069417E-01 .990305472E-05    3
-.119062354E-07 .290135824E-11-.249124705E+05 .642168604E+01                   4
C3H6O2                  C   3H   6O   2     G    300.00   4000.00 1382.00      1
 .118936666E+02 .144153203E-01-.477525443E-05 .726036430E-09-.415285995E-13    2
-.459271652E+05-.327285750E+02 .266613285E+01 .346302298E-01-.214380719E-04    3
 .690469334E-08-.916939105E-12-.425706030E+05 .173358364E+02                   4
ACETOL                  C   3H   6O   2     G    300.00   4000.00 1390.00      1
 .110277409E+02 .156022896E-01-.518498789E-05 .789604263E-09-.452017356E-13    2
-.493518932E+05-.296460029E+02 .170110573E+01 .349995386E-01-.195672111E-04    3
 .513929120E-08-.454830190E-12-.458857790E+05 .212715964E+02                   4
C3H5OOH                 C   3H   6O   2     G    300.00   4000.00 1382.00      1
 .139268456E+02 .135384067E-01-.474335693E-05 .748389157E-09-.439105886E-13    2
-.132537727E+05-.456757848E+02 .221491505E+01 .390935107E-01-.258809564E-04    3
 .870894601E-08-.120793929E-11-.896037969E+04 .179425329E+02                   4
C3-OQOOH                C   3H   6O   3     G    300.00   4000.00 1391.00      1
 .170285271E+02 .130716784E-01-.459310856E-05 .726135156E-09-.426658337E-13    2
-.416334217E+05-.592513577E+02 .768933034E+00 .546905880E-01-.465072405E-04    3
 .203159585E-07-.358398999E-11-.363238861E+05 .268291637E+02                   4
C3H8                    C   3H   8          G    300.00   4000.00 1000.00      1
 .752530602E+01 .188903400E-01-.628392400E-05 .917937280E-09-.481240960E-13    2
-.164646226E+05-.178445202E+02 .896921000E+00 .266898590E-01 .543142510E-05    3
-.212600000E-07 .924333010E-11-.139549200E+05 .193553300E+02                   4
NC3H7OH                 C   3H   8O   1     G    300.00   4000.00 1396.00      1
 .107520626E+02 .180260472E-01-.603049401E-05 .922166246E-09-.529319319E-13    2
-.361555719E+05-.310977038E+02 .978207214E-01 .420500918E-01-.267066894E-04    3
 .903941170E-08-.128324751E-11-.323437836E+05 .264700804E+02                   4
IC3H7OH                 C   3H   8O   1     G    300.00   4000.00 1000.00      1
 .577239007E+01 .268947430E-01-.111795290E-04 .211392460E-08-.149320990E-12    2
-.361710675E+05-.384089810E+01-.176838920E+00 .452559560E-01-.319190720E-04    3
 .123062880E-07-.201412540E-11-.346643940E+05 .263322250E+02                   4
C3H7OOH                 C   3H   8O   2     G    300.00   4000.00 1388.00      1
 .150655849E+02 .170865595E-01-.593183927E-05 .930136673E-09-.543384935E-13    2
-.301371140E+05-.515057998E+02 .783525746E+00 .504826223E-01-.365089942E-04    3
 .140377750E-07-.226737156E-11-.251105573E+05 .253041175E+02                   4
C4H2                    C   4H   2          G    300.00   4000.00 1000.00      1
 .903147468E+01 .604725210E-02-.194878790E-05 .275486300E-09-.138560800E-13    2
 .529472934E+05-.238511290E+02 .400519100E+01 .198100000E-01-.986587660E-05    3
-.663515820E-08 .607741290E-11 .542406400E+05 .184573600E+01                   4
C4H4                    C   4H   4          G    300.00   4000.00 1000.00      1
 .665080310E+01 .161294300E-01-.719388700E-05 .149817800E-08-.118641100E-12    2
 .311958636E+05-.979559836E+01-.191524700E+01 .527508700E-01-.716559400E-04    3
 .550724200E-07-.172862200E-10 .329785000E+05 .314199800E+02                   4
C4H6                    C   4H   6          G    300.00   4000.00 1000.00      1
 .823794980E+01 .173695890E-01-.615923200E-05 .979908060E-09-.578075590E-13    2
 .923259930E+04-.203418190E+02 .112443850E+00 .343711770E-01-.111106630E-04    3
-.921096660E-08 .620841700E-11 .118022620E+05 .230917180E+02                   4
C4H6O2                  C   4H   6O   2     G    300.00   4000.00 1375.00      1
 .135393551E+02 .168328392E-01-.587873230E-05 .925553795E-09-.542254877E-13    2
-.462482008E+05-.437360830E+02 .182538964E+01 .377978336E-01-.172044878E-04    3
 .195698878E-08 .398612932E-12-.415126261E+05 .214925508E+02                   4
IC4H8                   C   4H   8          G    300.00   4000.00 1388.00      1
 .112258330E+02 .181795798E-01-.620348592E-05 .961444458E-09-.557088057E-13    2
-.769983777E+04-.373306704E+02 .938433173E+00 .390547287E-01-.216437148E-04    3
 .587267077E-08-.614435479E-12-.374817891E+04 .191442985E+02                   4
NC4H8                   C   4H   8          G    300.00   4000.00 1000.00      1
 .205358410E+01 .343505070E-01-.158831970E-04 .330896620E-08-.253610450E-12    2
-.213972310E+04 .155432010E+02 .118113800E+01 .308533800E-01 .508652470E-05    3
-.246548880E-07 .111101930E-10-.179040040E+04 .210624690E+02                   4
CYC5H4O                 C   5H   4O   1     G    300.00   4000.00 1000.00      1
 .558734350E+01 .254149730E-01-.929145880E-05 .112347330E-08 .000000000E+00    2
 .339172461E+04-.552979995E+01-.427809100E+01 .546170700E-01-.380993520E-04    3
 .105947040E-07 .000000000E+00 .589093400E+04 .446629800E+02                   4
CYC5H6                  C   5H   6          G    300.00   4000.00 1000.00      1
 .230537462E+00 .409571826E-01-.241588958E-04 .679763480E-08-.736374421E-12    2
 .143779465E+05 .202551234E+02-.513691194E+01 .606953453E-01-.460552837E-04    3
 .128457201E-07 .741214852E-12 .153675713E+05 .461567559E+02                   4
C6H6                    C   6H   6          G    300.00   4000.00 1000.00      1
 .129109067E+02 .172329600E-01-.502421020E-05 .589349680E-09-.194752100E-13    2
 .366437279E+04-.500281184E+02-.313801200E+01 .472310300E-01-.296220700E-05    3
-.326281900E-07 .171869100E-10 .889003000E+04 .365757300E+02                   4
MCPTD                   C   6H   8          G    300.00   4000.00 1399.00      1
 .154352848E+02 .199801707E-01-.680270423E-05 .105349633E-08-.610336727E-13    2
 .447456576E+04-.636393642E+02-.665320026E+01 .744640477E-01-.582864186E-04    3
 .231603543E-07-.369017129E-11 .117669311E+05 .538162769E+02                   4
C10H8                   C  10H   8          G    300.00   4000.00 1401.00      1
 .234023214E+02 .242434427E-01-.836282016E-05 .130620111E-08-.761153748E-13    2
 .651941329E+04-.107433208E+03-.883645988E+01 .109300567E+00-.955200914E-04    3
 .421647669E-07-.739851710E-11 .166533366E+05 .621064766E+02                   4
N                       N   1               G    300.00   4000.00 1000.00      1
 .245026778E+01 .106614600E-03-.746533710E-07 .187965200E-10-.102598400E-14    2
 .561160257E+05 .444874779E+01 .250307100E+01-.218001810E-04 .542052910E-07    3
-.564755990E-10 .209990390E-13 .560988900E+05 .416756600E+01                   4
O                       O   1               G    300.00   4000.00 1000.00      1
 .254205876E+01-.275506100E-04-.310280290E-08 .455106700E-11-.436805100E-15    2
 .292307989E+05 .492030884E+01 .294642800E+01-.163816600E-02 .242103100E-05    3
-.160284300E-08 .389069610E-12 .291476400E+05 .296399500E+01                   4
NO3                     O   3N   1          G    300.00   4000.00 1000.00      1
 .712030587E+01 .324622800E-02-.143161340E-05 .279705300E-09-.201300700E-13    2
 .586448126E+04-.121372920E+02 .122107630E+01 .187879700E-01-.134432120E-04    3
 .127460130E-08 .135406010E-11 .747314400E+04 .184020200E+02                   4
H                       H   1               G    300.00   4000.00 1000.00      1
 .250000000E+01 .000000000E+00 .000000000E+00 .000000000E+00 .000000000E+00    2
 .254716200E+05-.460117600E+00 .250000000E+01 .000000000E+00 .000000000E+00    3
 .000000000E+00 .000000000E+00 .254716200E+05-.460117600E+00                   4
NH                      H   1N   1          G    300.00   4000.00 1000.00      1
 .276025108E+01 .137534600E-02-.445191400E-06 .769279080E-10-.501759190E-14    2
 .420782748E+05 .585718609E+01 .333975800E+01 .125300900E-02-.349164500E-05    3
 .421881200E-08-.155761800E-11 .418504700E+05 .250718000E+01                   4
NNH                     H   1N   2          G    300.00   4000.00 1000.00      1
 .441534072E+01 .161438800E-02-.163289400E-06-.855984590E-10 .161479110E-13    2
 .278802961E+05 .904297112E+00 .350134400E+01 .205358610E-02 .717040900E-06    3
 .492134780E-09-.967117010E-12 .283334700E+05 .639183800E+01                   4
OH                      H   1O   1          G    300.00   4000.00 1710.00      1
 .285376040E+01 .102994334E-02-.232666477E-06 .193750704E-10-.315759847E-15    2
 .369949720E+04 .578756825E+01 .341896226E+01 .319255801E-03-.308292717E-06    3
 .364407494E-09-.100195479E-12 .345264448E+04 .254433372E+01                   4
HO2                     H   1O   2          G    300.00   4000.00 1000.00      1
 .401721090E+01 .223982013E-02-.633658150E-06 .114246370E-09-.107908535E-13    2
 .111856713E+03 .378510215E+01 .430179801E+01-.474912051E-02 .211582891E-04    3
-.242763894E-07 .929225124E-11 .294808040E+03 .371666245E+01                   4
NH2                     H   2N   1          G    300.00   4000.00 1000.00      1
 .296131091E+01 .293269890E-02-.906360010E-06 .161725700E-09-.120420000E-13    2
 .219197637E+05 .577788090E+01 .343249300E+01 .329953990E-02-.661359990E-05    3
 .859094660E-08-.357204610E-11 .217722700E+05 .309011000E+01                   4
H2NO                    H   2O   1N   1     G    300.00   4000.00 1000.00      1
 .149675000E+01 .889472000E-02-.330837000E-05 .405760000E-09 .000000000E+00    2
 .724825208E+04 .175864616E+02 .267141000E+01 .529823000E-02 .360637000E-06    3
-.841417000E-09 .000000000E+00 .696062900E+04 .116499100E+02                   4
N2H3                    H   3N   2          G    300.00   4000.00 1000.00      1
 .444184100E+01 .721427100E-02-.249568400E-05 .392056500E-09-.229895000E-13    2
 .166422164E+05-.427486304E+00 .317420400E+01 .471590700E-02 .133486700E-04    3
-.191968500E-07 .748756400E-11 .172727000E+05 .755722400E+01                   4
C                       C   1               G    300.00   4000.00 1000.00      1
 .249266888E+01 .479889284E-04-.724335020E-07 .374291029E-10-.487277893E-14    2
 .854512953E+05 .480150373E+01 .255423955E+01-.321537724E-03 .733792245E-06    3
-.732234889E-09 .266521446E-12 .854438832E+05 .453130848E+01                   4
CN                      C   1N   1          G    300.00   4000.00 1000.00      1
 .372011754E+01 .151835110E-03 .198738110E-06-.379837100E-10 .132823000E-14    2
 .511162563E+05 .288861031E+01 .366320400E+01-.115652890E-02 .216340890E-05    3
 .185420800E-09-.821469520E-12 .512811700E+05 .373901500E+01                   4
NCN                     C   1N   2          G    300.00   4000.00 1000.00      1
 .568743460E+01 .182663439E-02-.707551130E-06 .119517763E-09-.731862017E-14    2
 .530454071E+05-.631950475E+01 .279807986E+01 .100008861E-01-.959242059E-05    3
 .475565678E-08-.104348512E-11 .538574577E+05 .862129570E+01                   4
NCO                     C   1O   1N   1     G    300.00   4000.00 1000.00      1
 .501204558E+01 .262677300E-02-.110824310E-05 .209385990E-09-.146034700E-13    2
 .173718555E+05-.183007911E+01 .283032000E+01 .887149010E-02-.894563620E-05    3
 .587691810E-08-.190773400E-11 .180054300E+05 .949883200E+01                   4
CH                      C   1H   1          G    300.00   4000.00 1000.00      1
 .219622115E+01 .234038100E-02-.705820130E-06 .900758220E-10-.385504010E-14    2
 .708672121E+05 .917838138E+01 .320020200E+01 .207287490E-02-.513443090E-05    3
 .573388980E-08-.195553300E-11 .704525700E+05 .333158700E+01                   4
HNCN                    C   1H   1N   2     G    300.00   4000.00 1000.00      1
 .553846448E+01 .389054126E-02-.138104752E-05 .221294765E-09-.131827325E-13    2
 .359635337E+05-.339587098E+01 .306754311E+01 .106789939E-01-.796224305E-05    3
 .259883390E-08-.127057612E-12 .366623508E+05 .941074995E+01                   4
HCO                     C   1H   1O   1     G    300.00   4000.00 1000.00      1
 .355727119E+01 .334557190E-02-.133500600E-05 .247057210E-09-.171385000E-13    2
 .391632208E+04 .555229973E+01 .289832900E+01 .619914620E-02-.962308420E-05    3
 .108982500E-07-.457488520E-11 .415992100E+04 .898361500E+01                   4
HCO3                    C   1H   1O   3     G    300.00   4000.00 1368.00      1
 .724073447E+01 .463312951E-02-.163693995E-05 .259706693E-09-.152964699E-13    2
-.187027386E+05-.649534993E+01 .396059309E+01 .106002279E-01-.525713351E-05    3
 .101716726E-08-.287487602E-13-.173599383E+05 .117807483E+02                   4
CH2S                    C   1H   2          G    300.00   4000.00 1000.00      1
 .355288641E+01 .206678800E-02-.191411600E-06-.110467300E-09 .202134890E-13    2
 .498497521E+05 .168658499E+01 .397126500E+01-.169908800E-03 .102536900E-05    3
 .249254990E-08-.198126610E-11 .498936700E+05 .575320760E-01                   4
CH2                     C   1H   2          G    300.00   4000.00 1000.00      1
 .363640757E+01 .193305600E-02-.168701600E-06-.100989900E-09 .180825510E-13    2
 .453413341E+05 .215656196E+01 .376223700E+01 .115981900E-02 .248958490E-06    3
 .880083620E-09-.733243490E-12 .453679000E+05 .171257700E+01                   4
H2CN                    C   1H   2N   1     G    300.00   4000.00 1000.00      1
 .520970151E+01 .296929110E-02-.285558910E-06-.163555000E-09 .304325890E-13    2
 .276771105E+05-.444446452E+01 .285166100E+01 .569523310E-02 .107114000E-05    3
-.162261200E-08-.235110810E-12 .286378200E+05 .899274900E+01                   4
CH3                     C   1H   3          G    300.00   4000.00 1000.00      1
 .284405718E+01 .613797410E-02-.223034500E-05 .378516110E-09-.245215900E-13    2
 .164378004E+05 .545265727E+01 .243044200E+01 .111241000E-01-.168022000E-04    3
 .162182910E-07-.586495220E-11 .164237800E+05 .678979400E+01                   4
CH2OH                   C   1H   3O   1     G    300.00   4000.00 1000.00      1
 .632751914E+01 .360827010E-02-.320154700E-06-.193875000E-09 .350970410E-13    2
-.447450931E+04-.832935988E+01 .286262800E+01 .100152700E-01-.528543520E-06    3
-.513853890E-08 .224604100E-11-.334967800E+04 .103979400E+02                   4
CH3O                    C   1H   3O   1     G    300.00   4000.00 1000.00      1
 .377081447E+01 .787149740E-02-.265638390E-05 .394443090E-09-.211261600E-13    2
 .127818951E+03 .292947482E+01 .210620400E+01 .721659510E-02 .533847200E-05    3
-.737763630E-08 .207561010E-11 .978601200E+03 .131521800E+02                   4
CH3OO                   C   1H   3O   2     G    300.00   4000.00 1385.00      1
 .595784570E+01 .790728626E-02-.268246234E-05 .413891337E-09-.239007330E-13    2
-.378178515E+03-.353671121E+01 .426146906E+01 .100873599E-01-.321506184E-05    3
 .209409267E-09 .418339103E-13 .473129653E+03 .634599067E+01                   4
C2N2                    C   2N   2          G    300.00   4000.00 1000.00      1
 .670549520E+01 .364271185E-02-.130939702E-05 .216421413E-09-.131193815E-13    2
 .348824335E+05-.104803146E+02 .232928126E+01 .261540993E-01-.490009889E-04    3
 .461923035E-07-.164325831E-10 .356900732E+05 .986348075E+01                   4
C2O                     C   2O   1          G    300.00   4000.00 1000.00      1
 .542468378E+01 .185393945E-02-.517932956E-06 .677646230E-10-.353315237E-14    2
 .437161379E+05-.369608405E+01 .286278214E+01 .119701204E-01-.180851222E-04    3
 .152777730E-07-.520063163E-11 .443125964E+05 .889759099E+01                   4
C2H                     C   2H   1          G    300.00   4000.00 1000.00      1
 .316780603E+01 .475221900E-02-.183787070E-05 .304190250E-09-.177232770E-13    2
 .671210651E+05 .663589763E+01 .288965730E+01 .134099610E-01-.284769500E-04    3
 .294791040E-07-.109331510E-10 .668393930E+05 .622296430E+01                   4
HCCO                    C   2H   1O   1     G    300.00   4000.00 1000.00      1
 .675807437E+01 .200040010E-02-.202760700E-06-.104113200E-09 .196516400E-13    2
 .190151261E+05-.907126528E+01 .504796600E+01 .445347790E-02 .226828210E-06    3
-.148209400E-08 .225074100E-12 .196589100E+05 .481843900E+00                   4
CH2CN                   C   2H   2N   1     G    300.00   4000.00 1000.00      1
 .460581482E+01 .944851600E-02-.471163290E-05 .113899570E-08-.108289420E-12    2
 .291714861E+05 .100843943E+01 .252967240E+01 .181141380E-01-.189605750E-04    3
 .119445830E-07-.325441420E-11 .295922930E+05 .109934410E+02                   4
C2H3                    C   2H   3          G    300.00   4000.00 1000.00      1
 .593346697E+01 .401774510E-02-.396673900E-06-.144126700E-09 .237864300E-13    2
 .318543468E+05-.853030497E+01 .245927600E+01 .737147590E-02 .210987200E-05    3
-.132164200E-08-.118478400E-11 .333522500E+05 .115562000E+02                   4
CH3CO                   C   2H   3O   1     G    300.00   4000.00 1000.00      1
 .561230883E+01 .844988600E-02-.285414690E-05 .423837600E-09-.226840300E-13    2
-.518788372E+04-.327515155E+01 .312527800E+01 .977822020E-02 .452144790E-05    3
-.900946160E-08 .319371700E-11-.410850700E+04 .112288500E+02                   4
CH2CHO                  C   2H   3O   1     G    300.00   4000.00 1500.00      1
 .971005743E+01 .385496600E-02-.467782500E-06-.150517900E-09 .294142800E-13    2
-.269248263E+04-.281056408E+02 .280220500E+00 .274031100E-01-.255468300E-04    3
 .130667900E-07-.275042500E-11 .668264800E+03 .223973100E+02                   4
CH3CO3                  C   2H   3O   3     G    300.00   4000.00 1000.00      1
 .102188027E+02 .888408630E-02-.222887620E-05 .166265570E-09 .000000000E+00    2
-.256023886E+05-.219354293E+02 .384065500E+01 .218595100E-01-.904528040E-05    3
 .385393800E-09 .000000000E+00-.234946000E+05 .124829900E+02                   4
C2H5                    C   2H   5          G    300.00   4000.00 1000.00      1
 .719047846E+01 .648407680E-02-.642806410E-06-.234787910E-09 .388087690E-13    2
 .106745471E+05-.147808755E+02 .269070100E+01 .871913320E-02 .441983820E-05    3
 .933870310E-09-.392777300E-11 .128704000E+05 .121382000E+02                   4
CH3CH2O                 C   2H   5O   1     G    300.00   4000.00 1389.00      1
 .787338637E+01 .113072907E-01-.384421421E-05 .594414105E-09-.343894538E-13    2
-.607273381E+04-.173415969E+02 .494420708E+00 .271774434E-01-.165909010E-04    3
 .515204200E-08-.648496915E-12-.335252925E+04 .228079378E+02                   4
CH3CHOH                 C   2H   5O   1     G    300.00   4000.00 1553.00      1
 .726570301E+01 .109588926E-01-.363662803E-05 .553659830E-09-.317012322E-13    2
-.864371441E+04-.106822851E+02 .183974631E+01 .187789371E-01-.460544253E-05    3
-.213116990E-08 .943772653E-12-.629595195E+04 .201446141E+02                   4
C2H4OH                  C   2H   5O   1     G    300.00   4000.00 1391.00      1
 .752244726E+01 .110492715E-01-.372576465E-05 .572827397E-09-.330061759E-13    2
-.729337464E+04-.124960750E+02 .117714711E+01 .248115685E-01-.150299503E-04    3
 .479006785E-08-.640994211E-12-.495369043E+04 .220081586E+02                   4
C2H5OO                  C   2H   5O   2     G    300.00   4000.00 1388.00      1
 .951115499E+01 .122676900E-01-.422364452E-05 .658474989E-09-.383095208E-13    2
-.676067578E+04-.223427083E+02 .177950508E+01 .304938087E-01-.216376209E-04    3
 .868906296E-08-.151788464E-11-.399101974E+04 .192919501E+02                   4
C2-QOOH                 C   2H   5O   2     G    300.00   4000.00 1396.00      1
 .116258666E+02 .100826346E-01-.347934362E-05 .543394220E-09-.316569294E-13    2
-.910568267E+03-.318522902E+02 .813237801E+00 .390063400E-01-.340643855E-04    3
 .155066226E-07-.284069840E-11 .250785787E+04 .249684459E+02                   4
C2-OOQOOH               C   2H   5O   4     G    300.00   4000.00 1387.00      1
 .145471032E+02 .123393823E-01-.427259469E-05 .668763337E-09-.390196721E-13    2
-.196338761E+05-.408784236E+02 .590031872E+01 .305658528E-01-.185905950E-04    3
 .567871605E-08-.702799577E-12-.163916571E+05 .633051038E+01                   4
C3H3                    C   3H   3          G    300.00   4000.00 1000.00      1
 .883104772E+01 .435719410E-02-.410906610E-06-.236872300E-09 .437652000E-13    2
 .384741917E+05-.217791939E+02 .475419900E+01 .110802800E-01 .279332310E-06    3
-.547921220E-08 .194962900E-11 .398888300E+05 .585454700E+00                   4
CH2CCH3                 C   3H   5          G    300.00   4000.00 1000.00      1
 .920976624E+01 .787141170E-02-.772452210E-06-.449735690E-09 .837727170E-13    2
 .285396699E+05-.223237088E+02 .316186300E+01 .151810000E-01 .272265900E-05    3
-.517711210E-08 .543528610E-13 .309554700E+05 .119797300E+02                   4
CH2CHCH2                C   3H   5          G    300.00   4000.00 1000.00      1
 .846871473E+01 .110576240E-01-.329817360E-05 .323385870E-09 .000000000E+00    2
 .160467269E+05-.206696057E+02 .227648600E+01 .198556410E-01 .112384200E-05    3
-.101457600E-07 .344134200E-11 .182949600E+05 .137251500E+02                   4
CHCHCH3                 C   3H   5          G    300.00   4000.00 1000.00      1
 .920976624E+01 .787141170E-02-.772452210E-06-.449735690E-09 .837727170E-13    2
 .285396699E+05-.223237088E+02 .316186300E+01 .151810000E-01 .272265900E-05    3
-.517711210E-08 .543528610E-13 .309554700E+05 .119797300E+02                   4
RALD3G                  C   3H   5O   1     G    300.00   4000.00 1375.00      1
 .870809249E+01 .169954492E-01-.678967812E-05 .115791412E-08-.713981613E-13    2
-.316945536E+04-.193250119E+02 .610490346E+01 .798359589E-02 .165150596E-04    3
-.148235750E-07 .341993565E-11-.416049715E+03 .575846684E+00                   4
CH3COCH2                C   3H   5O   1     G    300.00   4000.00 1391.00      1
 .102303674E+02 .116494161E-01-.401005537E-05 .625205246E-09-.363784362E-13    2
-.844376284E+04-.279195044E+02 .180339187E+01 .301407085E-01-.193505552E-04    3
 .638199034E-08-.866103180E-12-.537233261E+04 .178046408E+02                   4
RALD3B                  C   3H   5O   1     G    300.00   4000.00 1366.00      1
 .979372730E+01 .168079281E-01-.684815970E-05 .118460585E-08-.738195109E-13    2
-.875662870E+04-.294639062E+02 .667614768E+01 .261082031E-02 .280410577E-04    3
-.226802600E-07 .516442572E-11-.510504908E+04-.439698728E+01                   4
C3H5OO                  C   3H   5O   2     G    300.00   4000.00 1375.00      1
 .120289627E+02 .126220050E-01-.443107280E-05 .699998849E-09-.411059161E-13    2
 .440592543E+04-.346276747E+02 .316765415E+01 .300862111E-01-.169786280E-04    3
 .462955698E-08-.501220245E-12 .789477349E+04 .142601307E+02                   4
NC3H7                   C   3H   7          G    300.00   4000.00 1000.00      1
 .722715260E+01 .172648710E-01-.588880490E-05 .669183600E-09 .000000000E+00    2
 .782835831E+04-.127978858E+02 .192253600E+01 .247892700E-01 .181024900E-05    3
-.178326490E-07 .858299630E-11 .971328300E+04 .164927100E+02                   4
IC3H7                   C   3H   7          G    300.00   4000.00 1000.00      1
 .736341098E+01 .171331520E-01-.582028000E-05 .658834320E-09 .000000000E+00    2
 .604684608E+04-.148406654E+02 .171329900E+01 .254261610E-01 .158080800E-05    3
-.182128610E-07 .882771030E-11 .803580600E+04 .162790100E+02                   4
NC3H7O                  C   3H   7O   1     G    300.00   4000.00 1390.00      1
 .107032043E+02 .160908541E-01-.548805425E-05 .850429828E-09-.492755368E-13    2
-.101405419E+05-.313058764E+02-.595838475E+00 .410450833E-01-.263340323E-04    3
 .872638287E-08-.119115039E-11-.604569631E+04 .299328965E+02                   4
NC3-QOOH                C   3H   7O   2     G    300.00   4000.00 1374.00      1
 .146139980E+02 .143723015E-01-.488635144E-05 .756519620E-09-.438364992E-13    2
-.646101457E+04-.457478245E+02 .191005011E+01 .411666833E-01-.251630217E-04    3
 .711856873E-08-.698838732E-12-.179305093E+04 .234514457E+02                   4
IC3-QOOH                C   3H   7O   2     G    300.00   4000.00 1399.00      1
 .155030898E+02 .139802008E-01-.481811216E-05 .751835399E-09-.437743118E-13    2
-.741643030E+04-.523911482E+02-.184042862E+00 .564670638E-01-.501611253E-04    3
 .230526863E-07-.423866481E-11-.252333896E+04 .298354826E+02                   4
IC3H7OO                 C   3H   7O   2     G    300.00   4000.00 1392.00      1
 .132610651E+02 .162501084E-01-.558631798E-05 .870057473E-09-.505849469E-13    2
-.131937089E+05-.421023499E+02 .103495454E+01 .469942369E-01-.366525520E-04    3
 .157084173E-07-.281956117E-11-.906344820E+04 .229566921E+02                   4
NC3H7OO                 C   3H   7O   2     G    300.00   4000.00 1388.00      1
 .127230991E+02 .167336808E-01-.575943184E-05 .897769493E-09-.522275065E-13    2
-.108816595E+05-.381965321E+02 .156301709E+01 .426192697E-01-.296615075E-04    3
 .114187326E-07-.189894471E-11-.688086375E+04 .219842933E+02                   4
NC3-OOQOOH              C   3H   7O   4     G    300.00   4000.00 1388.00      1
 .185146106E+02 .164157074E-01-.573085844E-05 .901975314E-09-.528299084E-13    2
-.231819444E+05-.618247164E+02 .254387733E+01 .570847379E-01-.472164204E-04    3
 .208289492E-07-.378162942E-11-.178600410E+05 .229447574E+02                   4
IC3-OOQOOH              C   3H   7O   4     G    300.00   4000.00 1391.00      1
 .191234208E+02 .158457151E-01-.552231946E-05 .868162288E-09-.508094203E-13    2
-.255253957E+05-.661419362E+02 .175906535E+01 .624712381E-01-.554930416E-04    3
 .257973727E-07-.483190839E-11-.200009572E+05 .251348546E+02                   4
C4H3                    C   4H   3          G    300.00   4000.00 1000.00      1
 .107527376E+02 .538115300E-02-.554963720E-06-.305226590E-09 .576173970E-13    2
 .612141980E+05-.297302533E+02 .415388100E+01 .172628700E-01-.238937390E-06    3
-.101870000E-07 .434050410E-11 .633807200E+05 .603650600E+01                   4
C4H5                    C   4H   5          G    300.00   4000.00 1000.00      1
 .128659744E+02 .794336940E-02-.862646570E-06-.465563500E-09 .895113110E-13    2
 .378355213E+05-.418250446E+02 .299524000E+01 .228845610E-01 .197547090E-05    3
-.114824500E-07 .319782310E-11 .414221800E+05 .128945400E+02                   4
CH2C3H5                 C   4H   7          G    300.00   4000.00 1000.00      1
 .664945270E+01 .226232110E-01-.806420670E-05 .954149200E-09 .000000000E+00    2
 .206794519E+05-.786429084E+01 .283048200E+00 .386777000E-01-.210739710E-04    3
 .427582900E-08 .000000000E+00 .225247800E+05 .254564400E+02                   4
SC4H7                   C   4H   7          G    300.00   4000.00 1000.00      1
 .714879043E+01 .219663880E-01-.774471300E-05 .907477370E-09 .000000000E+00    2
 .124589843E+05-.117547735E+02-.442598200E+00 .422160100E-01-.254697900E-04    3
 .597432100E-08 .000000000E+00 .145672100E+05 .276086500E+02                   4
IC4H7                   C   4H   7          G    300.00   4000.00 1000.00      1
 .616543300E+01 .257842760E-01-.936521250E-05 .112618500E-08 .000000000E+00    2
 .114713700E+05-.676561500E+01 .476952000E+01 .167724920E-01 .213011010E-04    3
-.275874430E-07 .845501100E-11 .126384700E+05 .401309300E+01                   4
NC4H9P                  C   4H   9          G    300.00   4000.00 1000.00      1
 .285927140E+01 .339093470E-01-.129634890E-04 .162487360E-08 .000000000E+00    2
 .644131902E+04 .136765387E+02 .361027200E+00 .446560900E-01-.269622400E-04    3
 .737512580E-08 .000000000E+00 .679487900E+04 .252696800E+02                   4
NC4H9S                  C   4H   9          G    300.00   4000.00 1000.00      1
 .182440000E+01 .354350280E-01-.136901980E-04 .172985780E-08 .000000000E+00    2
 .521137543E+04 .190721830E+02 .882678800E+00 .419813690E-01-.239577090E-04    3
 .639274900E-08 .000000000E+00 .513670700E+04 .226104800E+02                   4
NC4H9-OO                C   4H   9O   2     G    300.00   4000.00 1392.00      1
 .164199470E+02 .207668293E-01-.714061871E-05 .111233445E-08-.646799300E-13    2
-.172909027E+05-.576444825E+02 .859225542E+00 .589774363E-01-.445935184E-04    3
 .184502497E-07-.321329944E-11-.119598721E+05 .254554544E+02                   4
CYC5H5                  C   5H   5          G    300.00   4000.00 1000.00      1
 .421464919E+01 .271834728E-01-.133173209E-04 .308980119E-08-.277879873E-12    2
 .288952416E+05-.305999781E-01-.737844042E+01 .972391818E-01-.169579138E-03    3
 .151818667E-06-.512075479E-10 .305514662E+05 .512829539E+02                   4
C5H5O                   C   5H   5O   1     G    300.00   4000.00 1395.00      1
 .149072105E+02 .136369619E-01-.470762207E-05 .736028654E-09-.429314124E-13    2
 .143724130E+05-.569296345E+02-.414628450E+01 .623584874E-01-.528374678E-04    3
 .224628793E-07-.380136191E-11 .204992627E+05 .437921058E+02                   4
NC5H9                   C   5H   9          G    300.00   4000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
C5EN-OO                 C   5H   9O   2     G    300.00   4000.00 1392.00      1
 .186695690E+02 .216228347E-01-.748565666E-05 .117148772E-08-.683420517E-13    2
-.458976288E+04-.678082548E+02 .338814185E+00 .676913346E-01-.538434525E-04    3
 .231725654E-07-.414643363E-11 .158489053E+04 .297116190E+02                   4
C6H5                    C   6H   5          G    300.00   4000.00 1000.00      1
 .157758892E+02 .965110900E-02-.942941600E-06-.546911100E-09 .102652200E-12    2
 .330269797E+05-.617628096E+02 .114355700E+00 .362732400E-01 .115828600E-05    3
-.219696400E-07 .846355600E-11 .383605400E+05 .238011700E+02                   4
